// ChaCha20 Decryption Module
// ChaCha20 is a symmetric stream cipher - decryption uses the same operation as encryption
// Decryption: ciphertext XOR keystream = plaintext
// The keystream is generated using the same quarter_round function and state matrix

module decryption #(
    parameter DATA_WIDTH = 32  // Can be configured for different data widths
)(
    input  logic [DATA_WIDTH-1:0] ciphertext,     // Encrypted data input
    input  logic [DATA_WIDTH-1:0] keystream,      // Keystream generated by ChaCha20 block function
    output logic [DATA_WIDTH-1:0] plaintext       // Decrypted data output
);

    // ChaCha20 decryption is simply XOR operation
    // Since encryption is: plaintext XOR keystream = ciphertext
    // Decryption is:       ciphertext XOR keystream = plaintext
    // This works because: (plaintext XOR keystream) XOR keystream = plaintext
    
    assign plaintext = ciphertext ^ keystream;

endmodule


// ChaCha20 Block Function Wrapper
// This generates the keystream used for both encryption and decryption
// Uses the quarter_round function internally (you'd need to build the full ChaCha20 block)

module chacha20_block (
    input  logic [31:0] key [8],           // 256-bit key (8 x 32-bit words)
    input  logic [31:0] nonce [3],         // 96-bit nonce (3 x 32-bit words)
    input  logic [31:0] counter,           // 32-bit block counter
    output logic [31:0] keystream [16]     // 512-bit keystream output (16 x 32-bit words)
);

    // ChaCha20 state matrix (16 words of 32 bits each)
    logic [31:0] state [16];
    logic [31:0] working_state [16];
    
    // Constants for ChaCha20 ("expand 32-byte k")
    localparam [31:0] CONST0 = 32'h61707865;  // "expa"
    localparam [31:0] CONST1 = 32'h3320646e;  // "nd 3"
    localparam [31:0] CONST2 = 32'h79622d32;  // "2-by"
    localparam [31:0] CONST3 = 32'h6b206574;  // "te k"

    // Initialize state matrix
    // Layout:
    // 0-3:   Constants
    // 4-11:  Key (256 bits)
    // 12:    Counter
    // 13-15: Nonce (96 bits)
    always_comb begin
        state[0]  = CONST0;
        state[1]  = CONST1;
        state[2]  = CONST2;
        state[3]  = CONST3;
        state[4]  = key[0];
        state[5]  = key[1];
        state[6]  = key[2];
        state[7]  = key[3];
        state[8]  = key[4];
        state[9]  = key[5];
        state[10] = key[6];
        state[11] = key[7];
        state[12] = counter;
        state[13] = nonce[0];
        state[14] = nonce[1];
        state[15] = nonce[2];
        
        // Copy to working state
        for (int i = 0; i < 16; i++) begin
            working_state[i] = state[i];
        end
        
        // NOTE: In a complete implementation, you would:
        // 1. Perform 20 rounds (10 double rounds) of quarter_round operations
        // 2. Each double round does:
        //    - Column rounds: QR on (0,4,8,12), (1,5,9,13), (2,6,10,14), (3,7,11,15)
        //    - Diagonal rounds: QR on (0,5,10,15), (1,6,11,12), (2,7,8,13), (3,4,9,14)
        // 3. Add the original state to the working state
        // 
        // For this example, we're showing the structure
        // In practice, you'd instantiate quarter_round modules here
        
        // Add original state to working state (final step)
        for (int i = 0; i < 16; i++) begin
            keystream[i] = working_state[i] + state[i];
        end
    end

endmodule


// Complete ChaCha20 Encryption/Decryption System
// Demonstrates the full encrypt/decrypt cycle

module chacha20_cipher #(
    parameter BLOCK_SIZE = 512  // ChaCha20 operates on 512-bit blocks
)(
    input  logic [31:0] key [8],           // 256-bit key
    input  logic [31:0] nonce [3],         // 96-bit nonce
    input  logic [31:0] counter,           // Block counter
    input  logic [31:0] data_in [16],      // Input data (plaintext or ciphertext)
    input  logic        mode,              // 0 = encrypt, 1 = decrypt (both do same thing!)
    output logic [31:0] data_out [16]      // Output data (ciphertext or plaintext)
);

    // Generate keystream
    logic [31:0] keystream [16];
    
    chacha20_block block_gen (
        .key(key),
        .nonce(nonce),
        .counter(counter),
        .keystream(keystream)
    );
    
    // XOR data with keystream (same operation for encrypt and decrypt!)
    genvar i;
    generate
        for (i = 0; i < 16; i++) begin : xor_loop
            decryption #(.DATA_WIDTH(32)) dec (
                .ciphertext(data_in[i]),
                .keystream(keystream[i]),
                .plaintext(data_out[i])
            );
        end
    endgenerate

endmodule
