// Luhn Algorithm Validator
// Validates a 16-digit decimal number using the Luhn algorithm
// Input: 16 digits (each 4 bits, BCD encoded)
// Output: valid (1 if checksum passes, 0 otherwise)

module luhn_validator (
    input  logic        pan_ready,
    input  logic [75:0] pan_bcd,   // digit0 at [3:0] (leftmost) ... digit15 at [63:60] (rightmost/check)
    output logic        valid
);

    // Internally keep the same digit convention:
    // digit[0] is rightmost (check digit), digit[15] is leftmost
    logic [3:0] digit [15:0];
    logic [3:0] processed [15:0];
    logic [8:0] total_sum;          // 9 bits are enough: max sum = 16*9 = 144 (< 2^9)

    integer i;

    always_comb begin
        // Map pan_bcd (leftmost-first) -> digit[] (rightmost-first)
        for (i = 0; i < 16; i = i + 1) begin
            digit[i] = pan_bcd[4*(15 - i) +: 4];
        end

        // Process digit 0 (rightmost) - no doubling
        processed[0] = digit[0];

        // Process digit 1 - double it
        if (digit[1] <= 4'd4) begin
            processed[1] = digit[1] << 1;  // Just double
        end else begin
            processed[1] = (digit[1] << 1) - 4'd9;  // Double and subtract 9 (adds digits)
        end

        // Process digit 2 - no doubling
        processed[2] = digit[2];

        // Process digit 3 - double it
        if (digit[3] <= 4'd4) begin
            processed[3] = digit[3] << 1;
        end else begin
            processed[3] = (digit[3] << 1) - 4'd9;
        end

        // Process digit 4 - no doubling
        processed[4] = digit[4];

        // Process digit 5 - double it
        if (digit[5] <= 4'd4) begin
            processed[5] = digit[5] << 1;
        end else begin
            processed[5] = (digit[5] << 1) - 4'd9;
        end

        // Process digit 6 - no doubling
        processed[6] = digit[6];

        // Process digit 7 - double it
        if (digit[7] <= 4'd4) begin
            processed[7] = digit[7] << 1;
        end else begin
            processed[7] = (digit[7] << 1) - 4'd9;
        end

        // Process digit 8 - no doubling
        processed[8] = digit[8];

        // Process digit 9 - double it
        if (digit[9] <= 4'd4) begin
            processed[9] = digit[9] << 1;
        end else begin
            processed[9] = (digit[9] << 1) - 4'd9;
        end

        // Process digit 10 - no doubling
        processed[10] = digit[10];

        // Process digit 11 - double it
        if (digit[11] <= 4'd4) begin
            processed[11] = digit[11] << 1;
        end else begin
            processed[11] = (digit[11] << 1) - 4'd9;
        end

        // Process digit 12 - no doubling
        processed[12] = digit[12];

        // Process digit 13 - double it
        if (digit[13] <= 4'd4) begin
            processed[13] = digit[13] << 1;
        end else begin
            processed[13] = (digit[13] << 1) - 4'd9;
        end

        // Process digit 14 - no doubling
        processed[14] = digit[14];

        // Process digit 15 - double it
        if (digit[15] <= 4'd4) begin
            processed[15] = digit[15] << 1;
        end else begin
            processed[15] = (digit[15] << 1) - 4'd9;
        end

        // ---------- FIXED SUM CALCULATION ----------
        total_sum = 9'd0;
        for (i = 0; i < 16; i = i + 1) begin
            // Zero‑extend each 4‑bit processed digit to 9 bits before adding
            total_sum = total_sum + {5'd0, processed[i]};
        end
        // -------------------------------------------

        // Valid if sum modulo 10 equals 0, and only meaningful once PAN capture is done
        valid = pan_ready && ((total_sum % 9'd10) == 9'd0);
    end

endmodule